//
// Disclaimer:
//
//   This Verilog source code is intended as a design reference
//   which illustrates how these types of functions can be implemented.
//   It is the user's responsibility to verify their design for
//   consistency and functionality through the use of formal
//   verification methods.  
//
// --------------------------------------------------------------------
//           
//                     Lih-Feng Tsaur
//                     UCSD CSE Department
//                     9500 Gilman Dr, La Jolla, CA 92093
//                     U.S.A
//
// --------------------------------------------------------------------
//
// Revision History : 0.0

module fulladder_tb;
reg a;
reg b;
reg c;
wire sum;
wire carry;

full_adder uut (  .a(a),   .b(b),.c(c),.sum(sum),.carry(carry)  );
initial begin
#10 a=1’b0;b=1’b0;c=1’b0;
#10 a=1’b0;b=1’b0;c=1’b1;
#10 a=1’b0;b=1’b1;c=1’b0;
#10 a=1’b0;b=1’b1;c=1’b1;
#10 a=1’b1;b=1’b0;c=1’b0;
#10 a=1’b1;b=1’b0;c=1’b1;
#10 a=1’b1;b=1’b1;c=1’b0;
#10 a=1’b1;b=1’b1;c=1’b1;
#10 $stop;
End

endmodule
